module model

[heap]
pub type Unit = struct {}

pub const unit = Unit{}
